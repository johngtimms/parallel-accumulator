// EE 454
// Spring 2015
// Lab 2 Part 2
// John Timms
// accumulator_top.v
//
// load wire is for testbench
//

`timescale 1 ns / 100 ps

module accumulator_top (bus_clk, proc_clk, reset, load, result);

input bus_clk, proc_clk, reset;
input [31:0] load;
output [31:0] result;

wire [3:0] req;
wire [3:0] grant;

wire [1:0] op;
wire [31:0] data;
wire load_signal, full;

assign load_signal = (load != 0) ? 1'b1 : 1'b0;
assign data = (load != 0) ? load : 32'bz;
assign result = (full) ? data : 32'b0;

RoundRobinArbiter 		arbiter	(bus_clk, req, grant);
accumulator_memory		memory	(proc_clk, reset, op, data, load_signal, full);
accumulator_processor 	proc0 	(proc_clk, reset, op, data, req[0], grant[0]);
accumulator_processor 	proc1 	(proc_clk, reset, op, data, req[1], grant[1]);
accumulator_processor	proc2 	(proc_clk, reset, op, data, req[2], grant[2]);
accumulator_processor 	proc3 	(proc_clk, reset, op, data, req[3], grant[3]);

endmodule
 